
module PCS_generator_tb;

  // Parameters
  localparam  DATA_WIDTH           = 64                                                                                                                                                                                                                                                     ;                          
  localparam  HDR_WIDTH            = 2                                                                                                                                                                                                                                                      ;                          
  localparam  FRAME_WIDTH          = DATA_WIDTH + HDR_WIDTH                                                                                                                                                                                                                                 ;                          
  localparam  CONTROL_WIDTH        = 8                                                                                                                                                                                                                                                      ;                          
  localparam  TRANSCODER_BLOCKS    = 4                                                                                                                                                                                                                                                      ;                                   
  localparam  TRANSCODER_WIDTH     = 257                                                                                                                                                                                                                                                    ;                              
  localparam  TRANSCODER_HDR_WIDTH = 4                                                                                                                                                                                                                                                      ;                          
  localparam  PROB                 = 30                                                                                                                                                                                                                                                     ;                          
              
  logic [TRANSCODER_WIDTH  - 1 : 0] o_tx_scrambled_f0   /* Output scrambler                       */                                                                                                                                                                                        ;
  logic [TRANSCODER_WIDTH  - 1 : 0] o_tx_scrambled_f1   /* Output scrambler                       */                                                                                                                                                                                        ;
  logic [TRANSCODER_WIDTH  - 1 : 0] o_tx_coded_f0       /* Output transcoder                      */                                                                                                                                                                                        ;
  logic [TRANSCODER_WIDTH  - 1 : 0] o_tx_coded_f1       /* Output transcoder                      */                                                                                                                                                                                        ;
  logic [FRAME_WIDTH       - 1 : 0] o_frame_0           /* Output frame 0                         */                                                                                                                                                                                        ;
  logic [FRAME_WIDTH       - 1 : 0] o_frame_1           /* Output frame 1                         */                                                                                                                                                                                        ;
  logic [FRAME_WIDTH       - 1 : 0] o_frame_2           /* Output frame 2                         */                                                                                                                                                                                        ;
  logic [FRAME_WIDTH       - 1 : 0] o_frame_3           /* Output frame 3                         */                                                                                                                                                                                        ;
  logic [FRAME_WIDTH       - 1 : 0] o_frame_4           /* Output frame 4                         */                                                                                                                                                                                        ;
  logic [FRAME_WIDTH       - 1 : 0] o_frame_5           /* Output frame 5                         */                                                                                                                                                                                        ;
  logic [FRAME_WIDTH       - 1 : 0] o_frame_6           /* Output frame 6                         */                                                                                                                                                                                        ;
  logic [FRAME_WIDTH       - 1 : 0] o_frame_7           /* Output frame 7                         */                                                                                                                                                                                        ;
  logic [DATA_WIDTH        - 1 : 0] i_txd               /* Input data                             */                                                                                                                                                                                        ;
  logic [CONTROL_WIDTH     - 1 : 0] i_txc               /* Input control byte                     */                                                                                                                                                                                        ;
  logic [TRANSCODER_BLOCKS - 1 : 0] i_data_sel_0        /* Data selector                          */                                                                                                                                                                                        ;
  logic [TRANSCODER_BLOCKS - 1 : 0] i_data_sel_1        /* Data selector                          */                                                                                                                                                                                        ;
  logic [2                     : 0] i_valid             /* Input to enable frame generation       */                                                                                                                                                                                        ;    
  logic                             i_enable            /* Flag to enable frame generation        */                                                                                                                                                                                        ;
  logic                             i_random_0          /* Flag to enable random frame generation */                                                                                                                                                                                        ;
  logic                             i_random_1          /* Flag to enable random frame generation */                                                                                                                                                                                        ;
  logic                             i_tx_test_mode      /* Flag to enable TX test mode            */                                                                                                                                                                                        ;
  logic                             i_rst_n             /* Reset                                  */                                                                                                                                                                                        ;    
  logic                             clk                 /* Clock                                  */                                                                                                                                                                                        ;      
              


  PCS_generator # (
    .DATA_WIDTH           (DATA_WIDTH           )                                                                                                                                                                                                                                           ,
    .HDR_WIDTH            (HDR_WIDTH            )                                                                                                                                                                                                                                           ,
    .FRAME_WIDTH          (FRAME_WIDTH          )                                                                                                                                                                                                                                           ,
    .CONTROL_WIDTH        (CONTROL_WIDTH        )                                                                                                                                                                                                                                           ,
    .TRANSCODER_BLOCKS    (TRANSCODER_BLOCKS    )                                                                                                                                                                                                                                           ,
    .TRANSCODER_WIDTH     (TRANSCODER_WIDTH     )                                                                                                                                                                                                                                           ,
    .TRANSCODER_HDR_WIDTH (TRANSCODER_HDR_WIDTH )                                                                                                                                                                                                                                           ,
    .PROB                 (PROB                 )
  )
  PCS_generator_inst (                                                                            
    .o_tx_scrambled_f0    (o_tx_scrambled_f0    )                                                                                                                                                                                                                                           ,                        
    .o_tx_scrambled_f1    (o_tx_scrambled_f1    )                                                                                                                                                                                                                                           ,                        
    .o_tx_coded_f0        (o_tx_coded_f0        )                                                                                                                                                                                                                                           ,                       
    .o_tx_coded_f1        (o_tx_coded_f1        )                                                                                                                                                                                                                                           ,               
    .o_frame_0            (o_frame_0            )                                                                                                                                                                                                                                           ,          
    .o_frame_1            (o_frame_1            )                                                                                                                                                                                                                                           ,                       
    .o_frame_2            (o_frame_2            )                                                                                                                                                                                                                                           ,                        
    .o_frame_3            (o_frame_3            )                                                                                                                                                                                                                                           ,          
    .o_frame_4            (o_frame_4            )                                                                                                                                                                                                                                           ,                       
    .o_frame_5            (o_frame_5            )                                                                                                                                                                                                                                           ,                        
    .o_frame_6            (o_frame_6            )                                                                                                                                                                                                                                           ,                                                                                                                                                                                                                                                                                  
    .o_frame_7            (o_frame_7            )                                                                                                                                                                                                                                           ,                                                                                                                                                                                                                                                                                  
    .i_txd                (i_txd                )                                                                                                                                                                                                                                           ,                      
    .i_txc                (i_txc                )                                                                                                                                                                                                                                           ,
    .i_data_sel_0         (i_data_sel_0         )                                                                                                                                                                                                                                           ,                      
    .i_data_sel_1         (i_data_sel_1         )                                                                                                                                                                                                                                           ,                      
    .i_valid              (i_valid              )                                                                                                                                                                                                                                           ,                          
    .i_enable             (i_enable             )                                                                                                                                                                                                                                           ,
    .i_random_0           (i_random_0           )                                                                                                                                                                                                                                           ,                       
    .i_random_1           (i_random_1           )                                                                                                                                                                                                                                           ,                       
    .i_tx_test_mode       (i_tx_test_mode       )                                                                                                                                                                                                                                           ,                       
    .i_rst_n              (i_rst_n              )                                                                                                                                                                                                                                           ,                           
    .clk                  (clk                  )                                                                                                                                                                                                                                           
      
  );

always #5  clk = ~clk                                                                                                                                                                                                                                                                       ; 

initial begin
    clk             = 'b0                                                                                                                                                                                                                                                                   ;
    i_rst_n         = 'b0                                                                                                                                                                                                                                                                   ;
    i_data_sel_0    = 'b0000                                                                                                                                                                                                                                                                ;
    i_data_sel_1    = 'b0000                                                                                                                                                                                                                                                                ;
    i_enable        = 'b0                                                                                                                                                                                                                                                                   ;      
    i_valid         = 'b000                                                                                                                                                                                                                                                                 ;
    i_tx_test_mode  = 'b0                                                                                                                                                                                                                                                                   ;
    i_random_0      = 'b0                                                                                                                                                                                                                                                                   ;
    i_random_1      = 'b0                                                                                                                                                                                                                                                                   ;
    i_txd           = 'b0                                                                                                                                                                                                                                                                   ;
    i_txc           = 'b0                                                                                                                                                                                                                                                                   ;
    #100                                                                                                                                                                                                                                                                                    ;
    i_rst_n         = 1'b1                                                                                                                                                                                                                                                                  ;
    i_enable        = 1'b1                                                                                                                                                                                                                                                                  ;
    i_valid         = 3'b111                                                                                                                                                                                                                                                                ;
    i_random_0      = 1'b1                                                                                                                                                                                                                                                                  ;
    #1000                                                                                                                                                                                                                                                                                   ;  
    i_random_0      = 1'b0                                                                                                                                                                                                                                                                  ;
    #100                                                                                                                                                                                                                                                                                    ;
    i_data_sel_0    = 4'b0001                                                                                                                                                                                                                                                               ;
    #100                                                                                                                                                                                                                                                                                    ;
    i_data_sel_0    = 4'b0010                                                                                                                                                                                                                                                               ;
    #100                                                                                                                                                                                                                                                                                    ;
    i_data_sel_0    = 4'b0011                                                                                                                                                                                                                                                               ;
    #100                                                                                                                                                                                                                                                                                    ;
    i_data_sel_0    = 4'b0100                                                                                                                                                                                                                                                               ;
    #100                                                                                                                                                                                                                                                                                    ;
    i_data_sel_0    = 4'b0101                                                                                                                                                                                                                                                               ;
    #100                                                                                                                                                                                                                                                                                    ;
    i_data_sel_0    = 4'b0110                                                                                                                                                                                                                                                               ;
    #100                                                                                                                                                                                                                                                                                    ;
    i_data_sel_0    = 4'b0111                                                                                                                                                                                                                                                               ;
    #100                                                                                                                                                                                                                                                                                    ;
    i_data_sel_0    = 4'b1000                                                                                                                                                                                                                                                               ;
    #100                                                                                                                                                                                                                                                                                    ;
    i_data_sel_0    = 4'b1001                                                                                                                                                                                                                                                               ;
    #100                                                                                                                                                                                                                                                                                    ;
    i_data_sel_0    = 4'b1010                                                                                                                                                                                                                                                               ;
    #100                                                                                                                                                                                                                                                                                    ;
    i_data_sel_0    = 4'b1011                                                                                                                                                                                                                                                               ;
    #100                                                                                                                                                                                                                                                                                    ;
    i_data_sel_0    = 4'b1100                                                                                                                                                                                                                                                               ;
    #100                                                                                                                                                                                                                                                                                    ;
    i_data_sel_0    = 4'b1101                                                                                                                                                                                                                                                               ;
    #100                                                                                                                                                                                                                                                                                    ;
    i_data_sel_0    = 4'b1110                                                                                                                                                                                                                                                               ;
    #100                                                                                                                                                                                                                                                                                    ;
    i_random_0      = 1'b1                                                                                                                                                                                                                                                                  ;
    #100                                                                                                                                                                                                                                                                                    ;
    i_valid         = 3'b000                                                                                                                                                                                                                                                                ; 
    #100                                                                                                                                                                                                                                                                                    ;
    i_valid         = 3'b001                                                                                                                                                                                                                                                                ;
    #100                                                                                                                                                                                                                                                                                    ;
    i_valid         = 3'b010                                                                                                                                                                                                                                                                ;
    #100                                                                                                                                                                                                                                                                                    ;
    i_valid         = 3'b011                                                                                                                                                                                                                                                                ;
    #100                                                                                                                                                                                                                                                                                    ;
    i_valid         = 3'b100                                                                                                                                                                                                                                                                ;
    #100                                                                                                                                                                                                                                                                                    ;
    i_valid         = 3'b101                                                                                                                                                                                                                                                                ;
    #100                                                                                                                                                                                                                                                                                    ;
    i_valid         = 3'b110                                                                                                                                                                                                                                                                ;
    #100                                                                                                                                                                                                                                                                                    ;
    i_valid         = 3'b111                                                                                                                                                                                                                                                                ;
    i_tx_test_mode  = 1'b1                                                                                                                                                                                                                                                                  ;
    #100                                                                                                                                                                                                                                                                                    ;
    i_tx_test_mode  = 1'b0                                                                                                                                                                                                                                                                  ;
    i_enable        = 1'b0                                                                                                                                                                                                                                                                  ;
    i_txc           = 8'h00                                                                                                                                                                                                                                                                 ;
    i_txd           = 64'hAAAAAAAAAAAAAAAA                                                                                                                                                                                                                                                  ;
    #10                                                                                                                                                                                                                                                                                     ;
    i_txd           = 64'h3333333333333333                                                                                                                                                                                                                                                  ;
    #10                                                                                                                                                                                                                                                                                     ;
    i_txd           = 64'h5555555555555555                                                                                                                                                                                                                                                  ;
    #10                                                                                                                                                                                                                                                                                     ;
    i_txd           = 64'hDDDDDDDDDDDDDDDD                                                                                                                                                                                                                                                  ;
    #10                                                                                                                                                                                                                                                                                     ;
    i_txd           = 64'h7777777777777777                                                                                                                                                                                                                                                  ;
    #10                                                                                                                                                                                                                                                                                     ;
    i_txd = 64'hFFFFFFFFFFFFFFFF                                                                                                                                                                                                                                                            ;
    #10                                                                                                                                                                                                                                                                                     ;
    i_txd = 64'h0000000000000000                                                                                                                                                                                                                                                            ;
    #10                                                                                                                                                                                                                                                                                     ;
    i_txd = 64'h1111111111111111                                                                                                                                                                                                                                                            ;
    #400                                                                                                                                                                                                                                                                                    ;
    $finish                                                                                                                                                                                                                                                                                 ;
end


endmodule