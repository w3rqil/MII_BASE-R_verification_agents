// Change to PRBS8 mode
i_pattern_mode = PRBS8;
